module xnor_gate(a,b,o);
 	input a,b;
	output o;
	xnor g1(o,a,b);
endmodule



