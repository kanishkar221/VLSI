module nor_gate(a,b,o);
input a,b;
output o;
nor g1(o,a,b);  
endmodule



