module xor_gate(a,b,o);
	input a,b;
	output o;
	xor g1(o,a,b);
endmodule


