module and_gate (output Y, input A, B);
    and g1 (Y, A, B);  
endmodule
