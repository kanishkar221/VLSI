module not_gate(a,o);
	input a;
	output o;
	not g1(o,a);
endmodule



